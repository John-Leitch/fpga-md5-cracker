library verilog;
use verilog.vl_types.all;
entity Md5CoreTest is
end Md5CoreTest;
