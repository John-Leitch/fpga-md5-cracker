module Md5Core (
  input wire clk, 
  input wire [511:0] wb, 
  input wire [31:0] a0,
  input wire [31:0] b0, 
  input wire [31:0] c0, 
  input wire [31:0] d0, 
  output reg [31:0] a64, 
  output reg [31:0] b64, 
  output reg [31:0] c64, 
  output reg [31:0] d64);
  
  wire [31:0] w0 [0:15];
  assign w0[0] = wb[31:0];
  assign w0[1] = wb[63:32];
  assign w0[2] = wb[95:64];
  assign w0[3] = wb[127:96];
  assign w0[4] = wb[159:128];
  assign w0[5] = wb[191:160];
  assign w0[6] = wb[223:192];
  assign w0[7] = wb[255:224];
  assign w0[8] = wb[287:256];
  assign w0[9] = wb[319:288];
  assign w0[10] = wb[351:320];
  assign w0[11] = wb[383:352];
  assign w0[12] = wb[415:384];
  assign w0[13] = wb[447:416];
  assign w0[14] = wb[479:448];
  assign w0[15] = wb[511:480];

  reg [31:0] 
  a1, b1, c1, d1,
a2, b2, c2, d2,
a3, b3, c3, d3,
a4, b4, c4, d4,
a5, b5, c5, d5,
a6, b6, c6, d6,
a7, b7, c7, d7,
a8, b8, c8, d8,
a9, b9, c9, d9,
a10, b10, c10, d10,
a11, b11, c11, d11,
a12, b12, c12, d12,
a13, b13, c13, d13,
a14, b14, c14, d14,
a15, b15, c15, d15,
a16, b16, c16, d16,
a17, b17, c17, d17,
a18, b18, c18, d18,
a19, b19, c19, d19,
a20, b20, c20, d20,
a21, b21, c21, d21,
a22, b22, c22, d22,
a23, b23, c23, d23,
a24, b24, c24, d24,
a25, b25, c25, d25,
a26, b26, c26, d26,
a27, b27, c27, d27,
a28, b28, c28, d28,
a29, b29, c29, d29,
a30, b30, c30, d30,
a31, b31, c31, d31,
a32, b32, c32, d32,
a33, b33, c33, d33,
a34, b34, c34, d34,
a35, b35, c35, d35,
a36, b36, c36, d36,
a37, b37, c37, d37,
a38, b38, c38, d38,
a39, b39, c39, d39,
a40, b40, c40, d40,
a41, b41, c41, d41,
a42, b42, c42, d42,
a43, b43, c43, d43,
a44, b44, c44, d44,
a45, b45, c45, d45,
a46, b46, c46, d46,
a47, b47, c47, d47,
a48, b48, c48, d48,
a49, b49, c49, d49,
a50, b50, c50, d50,
a51, b51, c51, d51,
a52, b52, c52, d52,
a53, b53, c53, d53,
a54, b54, c54, d54,
a55, b55, c55, d55,
a56, b56, c56, d56,
a57, b57, c57, d57,
a58, b58, c58, d58,
a59, b59, c59, d59,
a60, b60, c60, d60,
a61, b61, c61, d61,
a62, b62, c62, d62,
a63, b63, c63, d63
; 

reg [31:0] w1 [0:15];
reg [31:0] w2 [0:15];
reg [31:0] w3 [0:15];
reg [31:0] w4 [0:15];
reg [31:0] w5 [0:15];
reg [31:0] w6 [0:15];
reg [31:0] w7 [0:15];
reg [31:0] w8 [0:15];
reg [31:0] w9 [0:15];
reg [31:0] w10 [0:15];
reg [31:0] w11 [0:15];
reg [31:0] w12 [0:15];
reg [31:0] w13 [0:15];
reg [31:0] w14 [0:15];
reg [31:0] w15 [0:15];
reg [31:0] w16 [0:15];
reg [31:0] w17 [0:15];
reg [31:0] w18 [0:15];
reg [31:0] w19 [0:15];
reg [31:0] w20 [0:15];
reg [31:0] w21 [0:15];
reg [31:0] w22 [0:15];
reg [31:0] w23 [0:15];
reg [31:0] w24 [0:15];
reg [31:0] w25 [0:15];
reg [31:0] w26 [0:15];
reg [31:0] w27 [0:15];
reg [31:0] w28 [0:15];
reg [31:0] w29 [0:15];
reg [31:0] w30 [0:15];
reg [31:0] w31 [0:15];
reg [31:0] w32 [0:15];
reg [31:0] w33 [0:15];
reg [31:0] w34 [0:15];
reg [31:0] w35 [0:15];
reg [31:0] w36 [0:15];
reg [31:0] w37 [0:15];
reg [31:0] w38 [0:15];
reg [31:0] w39 [0:15];
reg [31:0] w40 [0:15];
reg [31:0] w41 [0:15];
reg [31:0] w42 [0:15];
reg [31:0] w43 [0:15];
reg [31:0] w44 [0:15];
reg [31:0] w45 [0:15];
reg [31:0] w46 [0:15];
reg [31:0] w47 [0:15];
reg [31:0] w48 [0:15];
reg [31:0] w49 [0:15];
reg [31:0] w50 [0:15];
reg [31:0] w51 [0:15];
reg [31:0] w52 [0:15];
reg [31:0] w53 [0:15];
reg [31:0] w54 [0:15];
reg [31:0] w55 [0:15];
reg [31:0] w56 [0:15];
reg [31:0] w57 [0:15];
reg [31:0] w58 [0:15];
reg [31:0] w59 [0:15];
reg [31:0] w60 [0:15];
reg [31:0] w61 [0:15];
reg [31:0] w62 [0:15];
reg [31:0] w63 [0:15];


  
  always @(posedge clk)
    begin

a1 <= d0;
d1 <= c0;
c1 <= b0;
b1 <= b0 + ((((a0 + ((b0 & c0) | ((~b0) & d0)) + 'hd76aa478 + w0[0]) << 7) | ((a0 + ((b0 & c0) | ((~b0) & d0)) + 'hd76aa478 + w0[0]) >> (32 - 7))));
w1[0] <= w0[0];
w1[1] <= w0[1];
w1[2] <= w0[2];
w1[3] <= w0[3];
w1[4] <= w0[4];
w1[5] <= w0[5];
w1[6] <= w0[6];
w1[7] <= w0[7];
w1[8] <= w0[8];
w1[9] <= w0[9];
w1[10] <= w0[10];
w1[11] <= w0[11];
w1[12] <= w0[12];
w1[13] <= w0[13];
w1[14] <= w0[14];
w1[15] <= w0[15];

a2 <= d1;
d2 <= c1;
c2 <= b1;
b2 <= b1 + (((a1 + ((b1 & c1) | ((~b1) & d1)) + 'he8c7b756 + w1[1]) << 12) | ((a1 + ((b1 & c1) | ((~b1) & d1)) + 'he8c7b756 + w1[1]) >> (32 - 12)));
w2[0] <= w1[0];
w2[1] <= w1[1];
w2[2] <= w1[2];
w2[3] <= w1[3];
w2[4] <= w1[4];
w2[5] <= w1[5];
w2[6] <= w1[6];
w2[7] <= w1[7];
w2[8] <= w1[8];
w2[9] <= w1[9];
w2[10] <= w1[10];
w2[11] <= w1[11];
w2[12] <= w1[12];
w2[13] <= w1[13];
w2[14] <= w1[14];
w2[15] <= w1[15];

a3 <= d2;
d3 <= c2;
c3 <= b2;
b3 <= b2 + (((a2 + ((b2 & c2) | ((~b2) & d2)) + 'h242070db + w2[2]) << 17) | ((a2 + ((b2 & c2) | ((~b2) & d2)) + 'h242070db + w2[2]) >> (32 - 17)));
w3[0] <= w2[0];
w3[1] <= w2[1];
w3[2] <= w2[2];
w3[3] <= w2[3];
w3[4] <= w2[4];
w3[5] <= w2[5];
w3[6] <= w2[6];
w3[7] <= w2[7];
w3[8] <= w2[8];
w3[9] <= w2[9];
w3[10] <= w2[10];
w3[11] <= w2[11];
w3[12] <= w2[12];
w3[13] <= w2[13];
w3[14] <= w2[14];
w3[15] <= w2[15];

a4 <= d3;
d4 <= c3;
c4 <= b3;
b4 <= b3 + (((a3 + ((b3 & c3) | ((~b3) & d3)) + 'hc1bdceee + w3[3]) << 22) | ((a3 + ((b3 & c3) | ((~b3) & d3)) + 'hc1bdceee + w3[3]) >> (32 - 22)));
w4[0] <= w3[0];
w4[1] <= w3[1];
w4[2] <= w3[2];
w4[3] <= w3[3];
w4[4] <= w3[4];
w4[5] <= w3[5];
w4[6] <= w3[6];
w4[7] <= w3[7];
w4[8] <= w3[8];
w4[9] <= w3[9];
w4[10] <= w3[10];
w4[11] <= w3[11];
w4[12] <= w3[12];
w4[13] <= w3[13];
w4[14] <= w3[14];
w4[15] <= w3[15];

a5 <= d4;
d5 <= c4;
c5 <= b4;
b5 <= b4 + (((a4 + ((b4 & c4) | ((~b4) & d4)) + 'hf57c0faf + w4[4]) << 7) | ((a4 + ((b4 & c4) | ((~b4) & d4)) + 'hf57c0faf + w4[4]) >> (32 - 7)));
w5[0] <= w4[0];
w5[1] <= w4[1];
w5[2] <= w4[2];
w5[3] <= w4[3];
w5[4] <= w4[4];
w5[5] <= w4[5];
w5[6] <= w4[6];
w5[7] <= w4[7];
w5[8] <= w4[8];
w5[9] <= w4[9];
w5[10] <= w4[10];
w5[11] <= w4[11];
w5[12] <= w4[12];
w5[13] <= w4[13];
w5[14] <= w4[14];
w5[15] <= w4[15];

a6 <= d5;
d6 <= c5;
c6 <= b5;
b6 <= b5 + (((a5 + ((b5 & c5) | ((~b5) & d5)) + 'h4787c62a + w5[5]) << 12) | ((a5 + ((b5 & c5) | ((~b5) & d5)) + 'h4787c62a + w5[5]) >> (32 - 12)));
w6[0] <= w5[0];
w6[1] <= w5[1];
w6[2] <= w5[2];
w6[3] <= w5[3];
w6[4] <= w5[4];
w6[5] <= w5[5];
w6[6] <= w5[6];
w6[7] <= w5[7];
w6[8] <= w5[8];
w6[9] <= w5[9];
w6[10] <= w5[10];
w6[11] <= w5[11];
w6[12] <= w5[12];
w6[13] <= w5[13];
w6[14] <= w5[14];
w6[15] <= w5[15];

a7 <= d6;
d7 <= c6;
c7 <= b6;
b7 <= b6 + (((a6 + ((b6 & c6) | ((~b6) & d6)) + 'ha8304613 + w6[6]) << 17) | ((a6 + ((b6 & c6) | ((~b6) & d6)) + 'ha8304613 + w6[6]) >> (32 - 17)));
w7[0] <= w6[0];
w7[1] <= w6[1];
w7[2] <= w6[2];
w7[3] <= w6[3];
w7[4] <= w6[4];
w7[5] <= w6[5];
w7[6] <= w6[6];
w7[7] <= w6[7];
w7[8] <= w6[8];
w7[9] <= w6[9];
w7[10] <= w6[10];
w7[11] <= w6[11];
w7[12] <= w6[12];
w7[13] <= w6[13];
w7[14] <= w6[14];
w7[15] <= w6[15];

a8 <= d7;
d8 <= c7;
c8 <= b7;
b8 <= b7 + (((a7 + ((b7 & c7) | ((~b7) & d7)) + 'hfd469501 + w7[7]) << 22) | ((a7 + ((b7 & c7) | ((~b7) & d7)) + 'hfd469501 + w7[7]) >> (32 - 22)));
w8[0] <= w7[0];
w8[1] <= w7[1];
w8[2] <= w7[2];
w8[3] <= w7[3];
w8[4] <= w7[4];
w8[5] <= w7[5];
w8[6] <= w7[6];
w8[7] <= w7[7];
w8[8] <= w7[8];
w8[9] <= w7[9];
w8[10] <= w7[10];
w8[11] <= w7[11];
w8[12] <= w7[12];
w8[13] <= w7[13];
w8[14] <= w7[14];
w8[15] <= w7[15];

a9 <= d8;
d9 <= c8;
c9 <= b8;
b9 <= b8 + (((a8 + ((b8 & c8) | ((~b8) & d8)) + 'h698098d8 + w8[8]) << 7) | ((a8 + ((b8 & c8) | ((~b8) & d8)) + 'h698098d8 + w8[8]) >> (32 - 7)));
w9[0] <= w8[0];
w9[1] <= w8[1];
w9[2] <= w8[2];
w9[3] <= w8[3];
w9[4] <= w8[4];
w9[5] <= w8[5];
w9[6] <= w8[6];
w9[7] <= w8[7];
w9[8] <= w8[8];
w9[9] <= w8[9];
w9[10] <= w8[10];
w9[11] <= w8[11];
w9[12] <= w8[12];
w9[13] <= w8[13];
w9[14] <= w8[14];
w9[15] <= w8[15];

a10 <= d9;
d10 <= c9;
c10 <= b9;
b10 <= b9 + (((a9 + ((b9 & c9) | ((~b9) & d9)) + 'h8b44f7af + w9[9]) << 12) | ((a9 + ((b9 & c9) | ((~b9) & d9)) + 'h8b44f7af + w9[9]) >> (32 - 12)));
w10[0] <= w9[0];
w10[1] <= w9[1];
w10[2] <= w9[2];
w10[3] <= w9[3];
w10[4] <= w9[4];
w10[5] <= w9[5];
w10[6] <= w9[6];
w10[7] <= w9[7];
w10[8] <= w9[8];
w10[9] <= w9[9];
w10[10] <= w9[10];
w10[11] <= w9[11];
w10[12] <= w9[12];
w10[13] <= w9[13];
w10[14] <= w9[14];
w10[15] <= w9[15];

a11 <= d10;
d11 <= c10;
c11 <= b10;
b11 <= b10 + (((a10 + ((b10 & c10) | ((~b10) & d10)) + 'hffff5bb1 + w10[10]) << 17) | ((a10 + ((b10 & c10) | ((~b10) & d10)) + 'hffff5bb1 + w10[10]) >> (32 - 17)));
w11[0] <= w10[0];
w11[1] <= w10[1];
w11[2] <= w10[2];
w11[3] <= w10[3];
w11[4] <= w10[4];
w11[5] <= w10[5];
w11[6] <= w10[6];
w11[7] <= w10[7];
w11[8] <= w10[8];
w11[9] <= w10[9];
w11[10] <= w10[10];
w11[11] <= w10[11];
w11[12] <= w10[12];
w11[13] <= w10[13];
w11[14] <= w10[14];
w11[15] <= w10[15];

a12 <= d11;
d12 <= c11;
c12 <= b11;
b12 <= b11 + (((a11 + ((b11 & c11) | ((~b11) & d11)) + 'h895cd7be + w11[11]) << 22) | ((a11 + ((b11 & c11) | ((~b11) & d11)) + 'h895cd7be + w11[11]) >> (32 - 22)));
w12[0] <= w11[0];
w12[1] <= w11[1];
w12[2] <= w11[2];
w12[3] <= w11[3];
w12[4] <= w11[4];
w12[5] <= w11[5];
w12[6] <= w11[6];
w12[7] <= w11[7];
w12[8] <= w11[8];
w12[9] <= w11[9];
w12[10] <= w11[10];
w12[11] <= w11[11];
w12[12] <= w11[12];
w12[13] <= w11[13];
w12[14] <= w11[14];
w12[15] <= w11[15];

a13 <= d12;
d13 <= c12;
c13 <= b12;
b13 <= b12 + (((a12 + ((b12 & c12) | ((~b12) & d12)) + 'h6b901122 + w12[12]) << 7) | ((a12 + ((b12 & c12) | ((~b12) & d12)) + 'h6b901122 + w12[12]) >> (32 - 7)));
w13[0] <= w12[0];
w13[1] <= w12[1];
w13[2] <= w12[2];
w13[3] <= w12[3];
w13[4] <= w12[4];
w13[5] <= w12[5];
w13[6] <= w12[6];
w13[7] <= w12[7];
w13[8] <= w12[8];
w13[9] <= w12[9];
w13[10] <= w12[10];
w13[11] <= w12[11];
w13[12] <= w12[12];
w13[13] <= w12[13];
w13[14] <= w12[14];
w13[15] <= w12[15];

a14 <= d13;
d14 <= c13;
c14 <= b13;
b14 <= b13 + (((a13 + ((b13 & c13) | ((~b13) & d13)) + 'hfd987193 + w13[13]) << 12) | ((a13 + ((b13 & c13) | ((~b13) & d13)) + 'hfd987193 + w13[13]) >> (32 - 12)));
w14[0] <= w13[0];
w14[1] <= w13[1];
w14[2] <= w13[2];
w14[3] <= w13[3];
w14[4] <= w13[4];
w14[5] <= w13[5];
w14[6] <= w13[6];
w14[7] <= w13[7];
w14[8] <= w13[8];
w14[9] <= w13[9];
w14[10] <= w13[10];
w14[11] <= w13[11];
w14[12] <= w13[12];
w14[13] <= w13[13];
w14[14] <= w13[14];
w14[15] <= w13[15];

a15 <= d14;
d15 <= c14;
c15 <= b14;
b15 <= b14 + (((a14 + ((b14 & c14) | ((~b14) & d14)) + 'ha679438e + w14[14]) << 17) | ((a14 + ((b14 & c14) | ((~b14) & d14)) + 'ha679438e + w14[14]) >> (32 - 17)));
w15[0] <= w14[0];
w15[1] <= w14[1];
w15[2] <= w14[2];
w15[3] <= w14[3];
w15[4] <= w14[4];
w15[5] <= w14[5];
w15[6] <= w14[6];
w15[7] <= w14[7];
w15[8] <= w14[8];
w15[9] <= w14[9];
w15[10] <= w14[10];
w15[11] <= w14[11];
w15[12] <= w14[12];
w15[13] <= w14[13];
w15[14] <= w14[14];
w15[15] <= w14[15];

a16 <= d15;
d16 <= c15;
c16 <= b15;
b16 <= b15 + (((a15 + ((b15 & c15) | ((~b15) & d15)) + 'h49b40821 + w15[15]) << 22) | ((a15 + ((b15 & c15) | ((~b15) & d15)) + 'h49b40821 + w15[15]) >> (32 - 22)));
w16[0] <= w15[0];
w16[1] <= w15[1];
w16[2] <= w15[2];
w16[3] <= w15[3];
w16[4] <= w15[4];
w16[5] <= w15[5];
w16[6] <= w15[6];
w16[7] <= w15[7];
w16[8] <= w15[8];
w16[9] <= w15[9];
w16[10] <= w15[10];
w16[11] <= w15[11];
w16[12] <= w15[12];
w16[13] <= w15[13];
w16[14] <= w15[14];
w16[15] <= w15[15];

a17 <= d16;
d17 <= c16;
c17 <= b16;
b17 <= b16 + (((a16 + ((d16 & b16) | ((~d16) & c16)) + 'hf61e2562 + w16[(5 * 16 + 1) % 16]) << 5) | ((a16 + ((d16 & b16) | ((~d16) & c16)) + 'hf61e2562 + w16[(5 * 16 + 1) % 16]) >> (32 - 5)));
w17[0] <= w16[0];
w17[1] <= w16[1];
w17[2] <= w16[2];
w17[3] <= w16[3];
w17[4] <= w16[4];
w17[5] <= w16[5];
w17[6] <= w16[6];
w17[7] <= w16[7];
w17[8] <= w16[8];
w17[9] <= w16[9];
w17[10] <= w16[10];
w17[11] <= w16[11];
w17[12] <= w16[12];
w17[13] <= w16[13];
w17[14] <= w16[14];
w17[15] <= w16[15];

a18 <= d17;
d18 <= c17;
c18 <= b17;
b18 <= b17 + (((a17 + ((d17 & b17) | ((~d17) & c17)) + 'hc040b340 + w17[(5 * 17 + 1) % 16]) << 9) | ((a17 + ((d17 & b17) | ((~d17) & c17)) + 'hc040b340 + w17[(5 * 17 + 1) % 16]) >> (32 - 9)));
w18[0] <= w17[0];
w18[1] <= w17[1];
w18[2] <= w17[2];
w18[3] <= w17[3];
w18[4] <= w17[4];
w18[5] <= w17[5];
w18[6] <= w17[6];
w18[7] <= w17[7];
w18[8] <= w17[8];
w18[9] <= w17[9];
w18[10] <= w17[10];
w18[11] <= w17[11];
w18[12] <= w17[12];
w18[13] <= w17[13];
w18[14] <= w17[14];
w18[15] <= w17[15];

a19 <= d18;
d19 <= c18;
c19 <= b18;
b19 <= b18 + (((a18 + ((d18 & b18) | ((~d18) & c18)) + 'h265e5a51 + w18[(5 * 18 + 1) % 16]) << 14) | ((a18 + ((d18 & b18) | ((~d18) & c18)) + 'h265e5a51 + w18[(5 * 18 + 1) % 16]) >> (32 - 14)));
w19[0] <= w18[0];
w19[1] <= w18[1];
w19[2] <= w18[2];
w19[3] <= w18[3];
w19[4] <= w18[4];
w19[5] <= w18[5];
w19[6] <= w18[6];
w19[7] <= w18[7];
w19[8] <= w18[8];
w19[9] <= w18[9];
w19[10] <= w18[10];
w19[11] <= w18[11];
w19[12] <= w18[12];
w19[13] <= w18[13];
w19[14] <= w18[14];
w19[15] <= w18[15];

a20 <= d19;
d20 <= c19;
c20 <= b19;
b20 <= b19 + (((a19 + ((d19 & b19) | ((~d19) & c19)) + 'he9b6c7aa + w19[(5 * 19 + 1) % 16]) << 20) | ((a19 + ((d19 & b19) | ((~d19) & c19)) + 'he9b6c7aa + w19[(5 * 19 + 1) % 16]) >> (32 - 20)));
w20[0] <= w19[0];
w20[1] <= w19[1];
w20[2] <= w19[2];
w20[3] <= w19[3];
w20[4] <= w19[4];
w20[5] <= w19[5];
w20[6] <= w19[6];
w20[7] <= w19[7];
w20[8] <= w19[8];
w20[9] <= w19[9];
w20[10] <= w19[10];
w20[11] <= w19[11];
w20[12] <= w19[12];
w20[13] <= w19[13];
w20[14] <= w19[14];
w20[15] <= w19[15];

a21 <= d20;
d21 <= c20;
c21 <= b20;
b21 <= b20 + (((a20 + ((d20 & b20) | ((~d20) & c20)) + 'hd62f105d + w20[(5 * 20 + 1) % 16]) << 5) | ((a20 + ((d20 & b20) | ((~d20) & c20)) + 'hd62f105d + w20[(5 * 20 + 1) % 16]) >> (32 - 5)));
w21[0] <= w20[0];
w21[1] <= w20[1];
w21[2] <= w20[2];
w21[3] <= w20[3];
w21[4] <= w20[4];
w21[5] <= w20[5];
w21[6] <= w20[6];
w21[7] <= w20[7];
w21[8] <= w20[8];
w21[9] <= w20[9];
w21[10] <= w20[10];
w21[11] <= w20[11];
w21[12] <= w20[12];
w21[13] <= w20[13];
w21[14] <= w20[14];
w21[15] <= w20[15];

a22 <= d21;
d22 <= c21;
c22 <= b21;
b22 <= b21 + (((a21 + ((d21 & b21) | ((~d21) & c21)) + 'h02441453 + w21[(5 * 21 + 1) % 16]) << 9) | ((a21 + ((d21 & b21) | ((~d21) & c21)) + 'h02441453 + w21[(5 * 21 + 1) % 16]) >> (32 - 9)));
w22[0] <= w21[0];
w22[1] <= w21[1];
w22[2] <= w21[2];
w22[3] <= w21[3];
w22[4] <= w21[4];
w22[5] <= w21[5];
w22[6] <= w21[6];
w22[7] <= w21[7];
w22[8] <= w21[8];
w22[9] <= w21[9];
w22[10] <= w21[10];
w22[11] <= w21[11];
w22[12] <= w21[12];
w22[13] <= w21[13];
w22[14] <= w21[14];
w22[15] <= w21[15];

a23 <= d22;
d23 <= c22;
c23 <= b22;
b23 <= b22 + (((a22 + ((d22 & b22) | ((~d22) & c22)) + 'hd8a1e681 + w22[(5 * 22 + 1) % 16]) << 14) | ((a22 + ((d22 & b22) | ((~d22) & c22)) + 'hd8a1e681 + w22[(5 * 22 + 1) % 16]) >> (32 - 14)));
w23[0] <= w22[0];
w23[1] <= w22[1];
w23[2] <= w22[2];
w23[3] <= w22[3];
w23[4] <= w22[4];
w23[5] <= w22[5];
w23[6] <= w22[6];
w23[7] <= w22[7];
w23[8] <= w22[8];
w23[9] <= w22[9];
w23[10] <= w22[10];
w23[11] <= w22[11];
w23[12] <= w22[12];
w23[13] <= w22[13];
w23[14] <= w22[14];
w23[15] <= w22[15];

a24 <= d23;
d24 <= c23;
c24 <= b23;
b24 <= b23 + (((a23 + ((d23 & b23) | ((~d23) & c23)) + 'he7d3fbc8 + w23[(5 * 23 + 1) % 16]) << 20) | ((a23 + ((d23 & b23) | ((~d23) & c23)) + 'he7d3fbc8 + w23[(5 * 23 + 1) % 16]) >> (32 - 20)));
w24[0] <= w23[0];
w24[1] <= w23[1];
w24[2] <= w23[2];
w24[3] <= w23[3];
w24[4] <= w23[4];
w24[5] <= w23[5];
w24[6] <= w23[6];
w24[7] <= w23[7];
w24[8] <= w23[8];
w24[9] <= w23[9];
w24[10] <= w23[10];
w24[11] <= w23[11];
w24[12] <= w23[12];
w24[13] <= w23[13];
w24[14] <= w23[14];
w24[15] <= w23[15];

a25 <= d24;
d25 <= c24;
c25 <= b24;
b25 <= b24 + (((a24 + ((d24 & b24) | ((~d24) & c24)) + 'h21e1cde6 + w24[(5 * 24 + 1) % 16]) << 5) | ((a24 + ((d24 & b24) | ((~d24) & c24)) + 'h21e1cde6 + w24[(5 * 24 + 1) % 16]) >> (32 - 5)));
w25[0] <= w24[0];
w25[1] <= w24[1];
w25[2] <= w24[2];
w25[3] <= w24[3];
w25[4] <= w24[4];
w25[5] <= w24[5];
w25[6] <= w24[6];
w25[7] <= w24[7];
w25[8] <= w24[8];
w25[9] <= w24[9];
w25[10] <= w24[10];
w25[11] <= w24[11];
w25[12] <= w24[12];
w25[13] <= w24[13];
w25[14] <= w24[14];
w25[15] <= w24[15];

a26 <= d25;
d26 <= c25;
c26 <= b25;
b26 <= b25 + (((a25 + ((d25 & b25) | ((~d25) & c25)) + 'hc33707d6 + w25[(5 * 25 + 1) % 16]) << 9) | ((a25 + ((d25 & b25) | ((~d25) & c25)) + 'hc33707d6 + w25[(5 * 25 + 1) % 16]) >> (32 - 9)));
w26[0] <= w25[0];
w26[1] <= w25[1];
w26[2] <= w25[2];
w26[3] <= w25[3];
w26[4] <= w25[4];
w26[5] <= w25[5];
w26[6] <= w25[6];
w26[7] <= w25[7];
w26[8] <= w25[8];
w26[9] <= w25[9];
w26[10] <= w25[10];
w26[11] <= w25[11];
w26[12] <= w25[12];
w26[13] <= w25[13];
w26[14] <= w25[14];
w26[15] <= w25[15];

a27 <= d26;
d27 <= c26;
c27 <= b26;
b27 <= b26 + (((a26 + ((d26 & b26) | ((~d26) & c26)) + 'hf4d50d87 + w26[(5 * 26 + 1) % 16]) << 14) | ((a26 + ((d26 & b26) | ((~d26) & c26)) + 'hf4d50d87 + w26[(5 * 26 + 1) % 16]) >> (32 - 14)));
w27[0] <= w26[0];
w27[1] <= w26[1];
w27[2] <= w26[2];
w27[3] <= w26[3];
w27[4] <= w26[4];
w27[5] <= w26[5];
w27[6] <= w26[6];
w27[7] <= w26[7];
w27[8] <= w26[8];
w27[9] <= w26[9];
w27[10] <= w26[10];
w27[11] <= w26[11];
w27[12] <= w26[12];
w27[13] <= w26[13];
w27[14] <= w26[14];
w27[15] <= w26[15];

a28 <= d27;
d28 <= c27;
c28 <= b27;
b28 <= b27 + (((a27 + ((d27 & b27) | ((~d27) & c27)) + 'h455a14ed + w27[(5 * 27 + 1) % 16]) << 20) | ((a27 + ((d27 & b27) | ((~d27) & c27)) + 'h455a14ed + w27[(5 * 27 + 1) % 16]) >> (32 - 20)));
w28[0] <= w27[0];
w28[1] <= w27[1];
w28[2] <= w27[2];
w28[3] <= w27[3];
w28[4] <= w27[4];
w28[5] <= w27[5];
w28[6] <= w27[6];
w28[7] <= w27[7];
w28[8] <= w27[8];
w28[9] <= w27[9];
w28[10] <= w27[10];
w28[11] <= w27[11];
w28[12] <= w27[12];
w28[13] <= w27[13];
w28[14] <= w27[14];
w28[15] <= w27[15];

a29 <= d28;
d29 <= c28;
c29 <= b28;
b29 <= b28 + (((a28 + ((d28 & b28) | ((~d28) & c28)) + 'ha9e3e905 + w28[(5 * 28 + 1) % 16]) << 5) | ((a28 + ((d28 & b28) | ((~d28) & c28)) + 'ha9e3e905 + w28[(5 * 28 + 1) % 16]) >> (32 - 5)));
w29[0] <= w28[0];
w29[1] <= w28[1];
w29[2] <= w28[2];
w29[3] <= w28[3];
w29[4] <= w28[4];
w29[5] <= w28[5];
w29[6] <= w28[6];
w29[7] <= w28[7];
w29[8] <= w28[8];
w29[9] <= w28[9];
w29[10] <= w28[10];
w29[11] <= w28[11];
w29[12] <= w28[12];
w29[13] <= w28[13];
w29[14] <= w28[14];
w29[15] <= w28[15];

a30 <= d29;
d30 <= c29;
c30 <= b29;
b30 <= b29 + (((a29 + ((d29 & b29) | ((~d29) & c29)) + 'hfcefa3f8 + w29[(5 * 29 + 1) % 16]) << 9) | ((a29 + ((d29 & b29) | ((~d29) & c29)) + 'hfcefa3f8 + w29[(5 * 29 + 1) % 16]) >> (32 - 9)));
w30[0] <= w29[0];
w30[1] <= w29[1];
w30[2] <= w29[2];
w30[3] <= w29[3];
w30[4] <= w29[4];
w30[5] <= w29[5];
w30[6] <= w29[6];
w30[7] <= w29[7];
w30[8] <= w29[8];
w30[9] <= w29[9];
w30[10] <= w29[10];
w30[11] <= w29[11];
w30[12] <= w29[12];
w30[13] <= w29[13];
w30[14] <= w29[14];
w30[15] <= w29[15];

a31 <= d30;
d31 <= c30;
c31 <= b30;
b31 <= b30 + (((a30 + ((d30 & b30) | ((~d30) & c30)) + 'h676f02d9 + w30[(5 * 30 + 1) % 16]) << 14) | ((a30 + ((d30 & b30) | ((~d30) & c30)) + 'h676f02d9 + w30[(5 * 30 + 1) % 16]) >> (32 - 14)));
w31[0] <= w30[0];
w31[1] <= w30[1];
w31[2] <= w30[2];
w31[3] <= w30[3];
w31[4] <= w30[4];
w31[5] <= w30[5];
w31[6] <= w30[6];
w31[7] <= w30[7];
w31[8] <= w30[8];
w31[9] <= w30[9];
w31[10] <= w30[10];
w31[11] <= w30[11];
w31[12] <= w30[12];
w31[13] <= w30[13];
w31[14] <= w30[14];
w31[15] <= w30[15];

a32 <= d31;
d32 <= c31;
c32 <= b31;
b32 <= b31 + (((a31 + ((d31 & b31) | ((~d31) & c31)) + 'h8d2a4c8a + w31[(5 * 31 + 1) % 16]) << 20) | ((a31 + ((d31 & b31) | ((~d31) & c31)) + 'h8d2a4c8a + w31[(5 * 31 + 1) % 16]) >> (32 - 20)));
w32[0] <= w31[0];
w32[1] <= w31[1];
w32[2] <= w31[2];
w32[3] <= w31[3];
w32[4] <= w31[4];
w32[5] <= w31[5];
w32[6] <= w31[6];
w32[7] <= w31[7];
w32[8] <= w31[8];
w32[9] <= w31[9];
w32[10] <= w31[10];
w32[11] <= w31[11];
w32[12] <= w31[12];
w32[13] <= w31[13];
w32[14] <= w31[14];
w32[15] <= w31[15];

a33 <= d32;
d33 <= c32;
c33 <= b32;
b33 <= b32 + (((a32 + (b32 ^ c32 ^ d32) + 'hfffa3942 + w32[(3 * 32 + 5) % 16]) << 4) | ((a32 + (b32 ^ c32 ^ d32) + 'hfffa3942 + w32[(3 * 32 + 5) % 16]) >> (32 - 4)));
w33[0] <= w32[0];
w33[1] <= w32[1];
w33[2] <= w32[2];
w33[3] <= w32[3];
w33[4] <= w32[4];
w33[5] <= w32[5];
w33[6] <= w32[6];
w33[7] <= w32[7];
w33[8] <= w32[8];
w33[9] <= w32[9];
w33[10] <= w32[10];
w33[11] <= w32[11];
w33[12] <= w32[12];
w33[13] <= w32[13];
w33[14] <= w32[14];
w33[15] <= w32[15];

a34 <= d33;
d34 <= c33;
c34 <= b33;
b34 <= b33 + (((a33 + (b33 ^ c33 ^ d33) + 'h8771f681 + w33[(3 * 33 + 5) % 16]) << 11) | ((a33 + (b33 ^ c33 ^ d33) + 'h8771f681 + w33[(3 * 33 + 5) % 16]) >> (32 - 11)));
w34[0] <= w33[0];
w34[1] <= w33[1];
w34[2] <= w33[2];
w34[3] <= w33[3];
w34[4] <= w33[4];
w34[5] <= w33[5];
w34[6] <= w33[6];
w34[7] <= w33[7];
w34[8] <= w33[8];
w34[9] <= w33[9];
w34[10] <= w33[10];
w34[11] <= w33[11];
w34[12] <= w33[12];
w34[13] <= w33[13];
w34[14] <= w33[14];
w34[15] <= w33[15];

a35 <= d34;
d35 <= c34;
c35 <= b34;
b35 <= b34 + (((a34 + (b34 ^ c34 ^ d34) + 'h6d9d6122 + w34[(3 * 34 + 5) % 16]) << 16) | ((a34 + (b34 ^ c34 ^ d34) + 'h6d9d6122 + w34[(3 * 34 + 5) % 16]) >> (32 - 16)));
w35[0] <= w34[0];
w35[1] <= w34[1];
w35[2] <= w34[2];
w35[3] <= w34[3];
w35[4] <= w34[4];
w35[5] <= w34[5];
w35[6] <= w34[6];
w35[7] <= w34[7];
w35[8] <= w34[8];
w35[9] <= w34[9];
w35[10] <= w34[10];
w35[11] <= w34[11];
w35[12] <= w34[12];
w35[13] <= w34[13];
w35[14] <= w34[14];
w35[15] <= w34[15];

a36 <= d35;
d36 <= c35;
c36 <= b35;
b36 <= b35 + (((a35 + (b35 ^ c35 ^ d35) + 'hfde5380c + w35[(3 * 35 + 5) % 16]) << 23) | ((a35 + (b35 ^ c35 ^ d35) + 'hfde5380c + w35[(3 * 35 + 5) % 16]) >> (32 - 23)));
w36[0] <= w35[0];
w36[1] <= w35[1];
w36[2] <= w35[2];
w36[3] <= w35[3];
w36[4] <= w35[4];
w36[5] <= w35[5];
w36[6] <= w35[6];
w36[7] <= w35[7];
w36[8] <= w35[8];
w36[9] <= w35[9];
w36[10] <= w35[10];
w36[11] <= w35[11];
w36[12] <= w35[12];
w36[13] <= w35[13];
w36[14] <= w35[14];
w36[15] <= w35[15];

a37 <= d36;
d37 <= c36;
c37 <= b36;
b37 <= b36 + (((a36 + (b36 ^ c36 ^ d36) + 'ha4beea44 + w36[(3 * 36 + 5) % 16]) << 4) | ((a36 + (b36 ^ c36 ^ d36) + 'ha4beea44 + w36[(3 * 36 + 5) % 16]) >> (32 - 4)));
w37[0] <= w36[0];
w37[1] <= w36[1];
w37[2] <= w36[2];
w37[3] <= w36[3];
w37[4] <= w36[4];
w37[5] <= w36[5];
w37[6] <= w36[6];
w37[7] <= w36[7];
w37[8] <= w36[8];
w37[9] <= w36[9];
w37[10] <= w36[10];
w37[11] <= w36[11];
w37[12] <= w36[12];
w37[13] <= w36[13];
w37[14] <= w36[14];
w37[15] <= w36[15];

a38 <= d37;
d38 <= c37;
c38 <= b37;
b38 <= b37 + (((a37 + (b37 ^ c37 ^ d37) + 'h4bdecfa9 + w37[(3 * 37 + 5) % 16]) << 11) | ((a37 + (b37 ^ c37 ^ d37) + 'h4bdecfa9 + w37[(3 * 37 + 5) % 16]) >> (32 - 11)));
w38[0] <= w37[0];
w38[1] <= w37[1];
w38[2] <= w37[2];
w38[3] <= w37[3];
w38[4] <= w37[4];
w38[5] <= w37[5];
w38[6] <= w37[6];
w38[7] <= w37[7];
w38[8] <= w37[8];
w38[9] <= w37[9];
w38[10] <= w37[10];
w38[11] <= w37[11];
w38[12] <= w37[12];
w38[13] <= w37[13];
w38[14] <= w37[14];
w38[15] <= w37[15];

a39 <= d38;
d39 <= c38;
c39 <= b38;
b39 <= b38 + (((a38 + (b38 ^ c38 ^ d38) + 'hf6bb4b60 + w38[(3 * 38 + 5) % 16]) << 16) | ((a38 + (b38 ^ c38 ^ d38) + 'hf6bb4b60 + w38[(3 * 38 + 5) % 16]) >> (32 - 16)));
w39[0] <= w38[0];
w39[1] <= w38[1];
w39[2] <= w38[2];
w39[3] <= w38[3];
w39[4] <= w38[4];
w39[5] <= w38[5];
w39[6] <= w38[6];
w39[7] <= w38[7];
w39[8] <= w38[8];
w39[9] <= w38[9];
w39[10] <= w38[10];
w39[11] <= w38[11];
w39[12] <= w38[12];
w39[13] <= w38[13];
w39[14] <= w38[14];
w39[15] <= w38[15];

a40 <= d39;
d40 <= c39;
c40 <= b39;
b40 <= b39 + (((a39 + (b39 ^ c39 ^ d39) + 'hbebfbc70 + w39[(3 * 39 + 5) % 16]) << 23) | ((a39 + (b39 ^ c39 ^ d39) + 'hbebfbc70 + w39[(3 * 39 + 5) % 16]) >> (32 - 23)));
w40[0] <= w39[0];
w40[1] <= w39[1];
w40[2] <= w39[2];
w40[3] <= w39[3];
w40[4] <= w39[4];
w40[5] <= w39[5];
w40[6] <= w39[6];
w40[7] <= w39[7];
w40[8] <= w39[8];
w40[9] <= w39[9];
w40[10] <= w39[10];
w40[11] <= w39[11];
w40[12] <= w39[12];
w40[13] <= w39[13];
w40[14] <= w39[14];
w40[15] <= w39[15];

a41 <= d40;
d41 <= c40;
c41 <= b40;
b41 <= b40 + (((a40 + (b40 ^ c40 ^ d40) + 'h289b7ec6 + w40[(3 * 40 + 5) % 16]) << 4) | ((a40 + (b40 ^ c40 ^ d40) + 'h289b7ec6 + w40[(3 * 40 + 5) % 16]) >> (32 - 4)));
w41[0] <= w40[0];
w41[1] <= w40[1];
w41[2] <= w40[2];
w41[3] <= w40[3];
w41[4] <= w40[4];
w41[5] <= w40[5];
w41[6] <= w40[6];
w41[7] <= w40[7];
w41[8] <= w40[8];
w41[9] <= w40[9];
w41[10] <= w40[10];
w41[11] <= w40[11];
w41[12] <= w40[12];
w41[13] <= w40[13];
w41[14] <= w40[14];
w41[15] <= w40[15];

a42 <= d41;
d42 <= c41;
c42 <= b41;
b42 <= b41 + (((a41 + (b41 ^ c41 ^ d41) + 'heaa127fa + w41[(3 * 41 + 5) % 16]) << 11) | ((a41 + (b41 ^ c41 ^ d41) + 'heaa127fa + w41[(3 * 41 + 5) % 16]) >> (32 - 11)));
w42[0] <= w41[0];
w42[1] <= w41[1];
w42[2] <= w41[2];
w42[3] <= w41[3];
w42[4] <= w41[4];
w42[5] <= w41[5];
w42[6] <= w41[6];
w42[7] <= w41[7];
w42[8] <= w41[8];
w42[9] <= w41[9];
w42[10] <= w41[10];
w42[11] <= w41[11];
w42[12] <= w41[12];
w42[13] <= w41[13];
w42[14] <= w41[14];
w42[15] <= w41[15];

a43 <= d42;
d43 <= c42;
c43 <= b42;
b43 <= b42 + (((a42 + (b42 ^ c42 ^ d42) + 'hd4ef3085 + w42[(3 * 42 + 5) % 16]) << 16) | ((a42 + (b42 ^ c42 ^ d42) + 'hd4ef3085 + w42[(3 * 42 + 5) % 16]) >> (32 - 16)));
w43[0] <= w42[0];
w43[1] <= w42[1];
w43[2] <= w42[2];
w43[3] <= w42[3];
w43[4] <= w42[4];
w43[5] <= w42[5];
w43[6] <= w42[6];
w43[7] <= w42[7];
w43[8] <= w42[8];
w43[9] <= w42[9];
w43[10] <= w42[10];
w43[11] <= w42[11];
w43[12] <= w42[12];
w43[13] <= w42[13];
w43[14] <= w42[14];
w43[15] <= w42[15];

a44 <= d43;
d44 <= c43;
c44 <= b43;
b44 <= b43 + (((a43 + (b43 ^ c43 ^ d43) + 'h04881d05 + w43[(3 * 43 + 5) % 16]) << 23) | ((a43 + (b43 ^ c43 ^ d43) + 'h04881d05 + w43[(3 * 43 + 5) % 16]) >> (32 - 23)));
w44[0] <= w43[0];
w44[1] <= w43[1];
w44[2] <= w43[2];
w44[3] <= w43[3];
w44[4] <= w43[4];
w44[5] <= w43[5];
w44[6] <= w43[6];
w44[7] <= w43[7];
w44[8] <= w43[8];
w44[9] <= w43[9];
w44[10] <= w43[10];
w44[11] <= w43[11];
w44[12] <= w43[12];
w44[13] <= w43[13];
w44[14] <= w43[14];
w44[15] <= w43[15];

a45 <= d44;
d45 <= c44;
c45 <= b44;
b45 <= b44 + (((a44 + (b44 ^ c44 ^ d44) + 'hd9d4d039 + w44[(3 * 44 + 5) % 16]) << 4) | ((a44 + (b44 ^ c44 ^ d44) + 'hd9d4d039 + w44[(3 * 44 + 5) % 16]) >> (32 - 4)));
w45[0] <= w44[0];
w45[1] <= w44[1];
w45[2] <= w44[2];
w45[3] <= w44[3];
w45[4] <= w44[4];
w45[5] <= w44[5];
w45[6] <= w44[6];
w45[7] <= w44[7];
w45[8] <= w44[8];
w45[9] <= w44[9];
w45[10] <= w44[10];
w45[11] <= w44[11];
w45[12] <= w44[12];
w45[13] <= w44[13];
w45[14] <= w44[14];
w45[15] <= w44[15];

a46 <= d45;
d46 <= c45;
c46 <= b45;
b46 <= b45 + (((a45 + (b45 ^ c45 ^ d45) + 'he6db99e5 + w45[(3 * 45 + 5) % 16]) << 11) | ((a45 + (b45 ^ c45 ^ d45) + 'he6db99e5 + w45[(3 * 45 + 5) % 16]) >> (32 - 11)));
w46[0] <= w45[0];
w46[1] <= w45[1];
w46[2] <= w45[2];
w46[3] <= w45[3];
w46[4] <= w45[4];
w46[5] <= w45[5];
w46[6] <= w45[6];
w46[7] <= w45[7];
w46[8] <= w45[8];
w46[9] <= w45[9];
w46[10] <= w45[10];
w46[11] <= w45[11];
w46[12] <= w45[12];
w46[13] <= w45[13];
w46[14] <= w45[14];
w46[15] <= w45[15];

a47 <= d46;
d47 <= c46;
c47 <= b46;
b47 <= b46 + (((a46 + (b46 ^ c46 ^ d46) + 'h1fa27cf8 + w46[(3 * 46 + 5) % 16]) << 16) | ((a46 + (b46 ^ c46 ^ d46) + 'h1fa27cf8 + w46[(3 * 46 + 5) % 16]) >> (32 - 16)));
w47[0] <= w46[0];
w47[1] <= w46[1];
w47[2] <= w46[2];
w47[3] <= w46[3];
w47[4] <= w46[4];
w47[5] <= w46[5];
w47[6] <= w46[6];
w47[7] <= w46[7];
w47[8] <= w46[8];
w47[9] <= w46[9];
w47[10] <= w46[10];
w47[11] <= w46[11];
w47[12] <= w46[12];
w47[13] <= w46[13];
w47[14] <= w46[14];
w47[15] <= w46[15];

a48 <= d47;
d48 <= c47;
c48 <= b47;
b48 <= b47 + (((a47 + (b47 ^ c47 ^ d47) + 'hc4ac5665 + w47[(3 * 47 + 5) % 16]) << 23) | ((a47 + (b47 ^ c47 ^ d47) + 'hc4ac5665 + w47[(3 * 47 + 5) % 16]) >> (32 - 23)));
w48[0] <= w47[0];
w48[1] <= w47[1];
w48[2] <= w47[2];
w48[3] <= w47[3];
w48[4] <= w47[4];
w48[5] <= w47[5];
w48[6] <= w47[6];
w48[7] <= w47[7];
w48[8] <= w47[8];
w48[9] <= w47[9];
w48[10] <= w47[10];
w48[11] <= w47[11];
w48[12] <= w47[12];
w48[13] <= w47[13];
w48[14] <= w47[14];
w48[15] <= w47[15];

a49 <= d48;
d49 <= c48;
c49 <= b48;
b49 <= b48 + (((a48 + (c48 ^ (b48 | (~d48))) + 'hf4292244 + w48[(7 * 48) % 16]) << 6) | ((a48 + (c48 ^ (b48 | (~d48))) + 'hf4292244 + w48[(7 * 48) % 16]) >> (32 - 6)));
w49[0] <= w48[0];
w49[1] <= w48[1];
w49[2] <= w48[2];
w49[3] <= w48[3];
w49[4] <= w48[4];
w49[5] <= w48[5];
w49[6] <= w48[6];
w49[7] <= w48[7];
w49[8] <= w48[8];
w49[9] <= w48[9];
w49[10] <= w48[10];
w49[11] <= w48[11];
w49[12] <= w48[12];
w49[13] <= w48[13];
w49[14] <= w48[14];
w49[15] <= w48[15];

a50 <= d49;
d50 <= c49;
c50 <= b49;
b50 <= b49 + (((a49 + (c49 ^ (b49 | (~d49))) + 'h432aff97 + w49[(7 * 49) % 16]) << 10) | ((a49 + (c49 ^ (b49 | (~d49))) + 'h432aff97 + w49[(7 * 49) % 16]) >> (32 - 10)));
w50[0] <= w49[0];
w50[1] <= w49[1];
w50[2] <= w49[2];
w50[3] <= w49[3];
w50[4] <= w49[4];
w50[5] <= w49[5];
w50[6] <= w49[6];
w50[7] <= w49[7];
w50[8] <= w49[8];
w50[9] <= w49[9];
w50[10] <= w49[10];
w50[11] <= w49[11];
w50[12] <= w49[12];
w50[13] <= w49[13];
w50[14] <= w49[14];
w50[15] <= w49[15];

a51 <= d50;
d51 <= c50;
c51 <= b50;
b51 <= b50 + (((a50 + (c50 ^ (b50 | (~d50))) + 'hab9423a7 + w50[(7 * 50) % 16]) << 15) | ((a50 + (c50 ^ (b50 | (~d50))) + 'hab9423a7 + w50[(7 * 50) % 16]) >> (32 - 15)));
w51[0] <= w50[0];
w51[1] <= w50[1];
w51[2] <= w50[2];
w51[3] <= w50[3];
w51[4] <= w50[4];
w51[5] <= w50[5];
w51[6] <= w50[6];
w51[7] <= w50[7];
w51[8] <= w50[8];
w51[9] <= w50[9];
w51[10] <= w50[10];
w51[11] <= w50[11];
w51[12] <= w50[12];
w51[13] <= w50[13];
w51[14] <= w50[14];
w51[15] <= w50[15];

a52 <= d51;
d52 <= c51;
c52 <= b51;
b52 <= b51 + (((a51 + (c51 ^ (b51 | (~d51))) + 'hfc93a039 + w51[(7 * 51) % 16]) << 21) | ((a51 + (c51 ^ (b51 | (~d51))) + 'hfc93a039 + w51[(7 * 51) % 16]) >> (32 - 21)));
w52[0] <= w51[0];
w52[1] <= w51[1];
w52[2] <= w51[2];
w52[3] <= w51[3];
w52[4] <= w51[4];
w52[5] <= w51[5];
w52[6] <= w51[6];
w52[7] <= w51[7];
w52[8] <= w51[8];
w52[9] <= w51[9];
w52[10] <= w51[10];
w52[11] <= w51[11];
w52[12] <= w51[12];
w52[13] <= w51[13];
w52[14] <= w51[14];
w52[15] <= w51[15];

a53 <= d52;
d53 <= c52;
c53 <= b52;
b53 <= b52 + (((a52 + (c52 ^ (b52 | (~d52))) + 'h655b59c3 + w52[(7 * 52) % 16]) << 6) | ((a52 + (c52 ^ (b52 | (~d52))) + 'h655b59c3 + w52[(7 * 52) % 16]) >> (32 - 6)));
w53[0] <= w52[0];
w53[1] <= w52[1];
w53[2] <= w52[2];
w53[3] <= w52[3];
w53[4] <= w52[4];
w53[5] <= w52[5];
w53[6] <= w52[6];
w53[7] <= w52[7];
w53[8] <= w52[8];
w53[9] <= w52[9];
w53[10] <= w52[10];
w53[11] <= w52[11];
w53[12] <= w52[12];
w53[13] <= w52[13];
w53[14] <= w52[14];
w53[15] <= w52[15];

a54 <= d53;
d54 <= c53;
c54 <= b53;
b54 <= b53 + (((a53 + (c53 ^ (b53 | (~d53))) + 'h8f0ccc92 + w53[(7 * 53) % 16]) << 10) | ((a53 + (c53 ^ (b53 | (~d53))) + 'h8f0ccc92 + w53[(7 * 53) % 16]) >> (32 - 10)));
w54[0] <= w53[0];
w54[1] <= w53[1];
w54[2] <= w53[2];
w54[3] <= w53[3];
w54[4] <= w53[4];
w54[5] <= w53[5];
w54[6] <= w53[6];
w54[7] <= w53[7];
w54[8] <= w53[8];
w54[9] <= w53[9];
w54[10] <= w53[10];
w54[11] <= w53[11];
w54[12] <= w53[12];
w54[13] <= w53[13];
w54[14] <= w53[14];
w54[15] <= w53[15];

a55 <= d54;
d55 <= c54;
c55 <= b54;
b55 <= b54 + (((a54 + (c54 ^ (b54 | (~d54))) + 'hffeff47d + w54[(7 * 54) % 16]) << 15) | ((a54 + (c54 ^ (b54 | (~d54))) + 'hffeff47d + w54[(7 * 54) % 16]) >> (32 - 15)));
w55[0] <= w54[0];
w55[1] <= w54[1];
w55[2] <= w54[2];
w55[3] <= w54[3];
w55[4] <= w54[4];
w55[5] <= w54[5];
w55[6] <= w54[6];
w55[7] <= w54[7];
w55[8] <= w54[8];
w55[9] <= w54[9];
w55[10] <= w54[10];
w55[11] <= w54[11];
w55[12] <= w54[12];
w55[13] <= w54[13];
w55[14] <= w54[14];
w55[15] <= w54[15];

a56 <= d55;
d56 <= c55;
c56 <= b55;
b56 <= b55 + (((a55 + (c55 ^ (b55 | (~d55))) + 'h85845dd1 + w55[(7 * 55) % 16]) << 21) | ((a55 + (c55 ^ (b55 | (~d55))) + 'h85845dd1 + w55[(7 * 55) % 16]) >> (32 - 21)));
w56[0] <= w55[0];
w56[1] <= w55[1];
w56[2] <= w55[2];
w56[3] <= w55[3];
w56[4] <= w55[4];
w56[5] <= w55[5];
w56[6] <= w55[6];
w56[7] <= w55[7];
w56[8] <= w55[8];
w56[9] <= w55[9];
w56[10] <= w55[10];
w56[11] <= w55[11];
w56[12] <= w55[12];
w56[13] <= w55[13];
w56[14] <= w55[14];
w56[15] <= w55[15];

a57 <= d56;
d57 <= c56;
c57 <= b56;
b57 <= b56 + (((a56 + (c56 ^ (b56 | (~d56))) + 'h6fa87e4f + w56[(7 * 56) % 16]) << 6) | ((a56 + (c56 ^ (b56 | (~d56))) + 'h6fa87e4f + w56[(7 * 56) % 16]) >> (32 - 6)));
w57[0] <= w56[0];
w57[1] <= w56[1];
w57[2] <= w56[2];
w57[3] <= w56[3];
w57[4] <= w56[4];
w57[5] <= w56[5];
w57[6] <= w56[6];
w57[7] <= w56[7];
w57[8] <= w56[8];
w57[9] <= w56[9];
w57[10] <= w56[10];
w57[11] <= w56[11];
w57[12] <= w56[12];
w57[13] <= w56[13];
w57[14] <= w56[14];
w57[15] <= w56[15];

a58 <= d57;
d58 <= c57;
c58 <= b57;
b58 <= b57 + (((a57 + (c57 ^ (b57 | (~d57))) + 'hfe2ce6e0 + w57[(7 * 57) % 16]) << 10) | ((a57 + (c57 ^ (b57 | (~d57))) + 'hfe2ce6e0 + w57[(7 * 57) % 16]) >> (32 - 10)));
w58[0] <= w57[0];
w58[1] <= w57[1];
w58[2] <= w57[2];
w58[3] <= w57[3];
w58[4] <= w57[4];
w58[5] <= w57[5];
w58[6] <= w57[6];
w58[7] <= w57[7];
w58[8] <= w57[8];
w58[9] <= w57[9];
w58[10] <= w57[10];
w58[11] <= w57[11];
w58[12] <= w57[12];
w58[13] <= w57[13];
w58[14] <= w57[14];
w58[15] <= w57[15];

a59 <= d58;
d59 <= c58;
c59 <= b58;
b59 <= b58 + (((a58 + (c58 ^ (b58 | (~d58))) + 'ha3014314 + w58[(7 * 58) % 16]) << 15) | ((a58 + (c58 ^ (b58 | (~d58))) + 'ha3014314 + w58[(7 * 58) % 16]) >> (32 - 15)));
w59[0] <= w58[0];
w59[1] <= w58[1];
w59[2] <= w58[2];
w59[3] <= w58[3];
w59[4] <= w58[4];
w59[5] <= w58[5];
w59[6] <= w58[6];
w59[7] <= w58[7];
w59[8] <= w58[8];
w59[9] <= w58[9];
w59[10] <= w58[10];
w59[11] <= w58[11];
w59[12] <= w58[12];
w59[13] <= w58[13];
w59[14] <= w58[14];
w59[15] <= w58[15];

a60 <= d59;
d60 <= c59;
c60 <= b59;
b60 <= b59 + (((a59 + (c59 ^ (b59 | (~d59))) + 'h4e0811a1 + w59[(7 * 59) % 16]) << 21) | ((a59 + (c59 ^ (b59 | (~d59))) + 'h4e0811a1 + w59[(7 * 59) % 16]) >> (32 - 21)));
w60[0] <= w59[0];
w60[1] <= w59[1];
w60[2] <= w59[2];
w60[3] <= w59[3];
w60[4] <= w59[4];
w60[5] <= w59[5];
w60[6] <= w59[6];
w60[7] <= w59[7];
w60[8] <= w59[8];
w60[9] <= w59[9];
w60[10] <= w59[10];
w60[11] <= w59[11];
w60[12] <= w59[12];
w60[13] <= w59[13];
w60[14] <= w59[14];
w60[15] <= w59[15];

a61 <= d60;
d61 <= c60;
c61 <= b60;
b61 <= b60 + (((a60 + (c60 ^ (b60 | (~d60))) + 'hf7537e82 + w60[(7 * 60) % 16]) << 6) | ((a60 + (c60 ^ (b60 | (~d60))) + 'hf7537e82 + w60[(7 * 60) % 16]) >> (32 - 6)));
w61[0] <= w60[0];
w61[1] <= w60[1];
w61[2] <= w60[2];
w61[3] <= w60[3];
w61[4] <= w60[4];
w61[5] <= w60[5];
w61[6] <= w60[6];
w61[7] <= w60[7];
w61[8] <= w60[8];
w61[9] <= w60[9];
w61[10] <= w60[10];
w61[11] <= w60[11];
w61[12] <= w60[12];
w61[13] <= w60[13];
w61[14] <= w60[14];
w61[15] <= w60[15];

a62 <= d61;
d62 <= c61;
c62 <= b61;
b62 <= b61 + (((a61 + (c61 ^ (b61 | (~d61))) + 'hbd3af235 + w61[(7 * 61) % 16]) << 10) | ((a61 + (c61 ^ (b61 | (~d61))) + 'hbd3af235 + w61[(7 * 61) % 16]) >> (32 - 10)));
w62[0] <= w61[0];
w62[1] <= w61[1];
w62[2] <= w61[2];
w62[3] <= w61[3];
w62[4] <= w61[4];
w62[5] <= w61[5];
w62[6] <= w61[6];
w62[7] <= w61[7];
w62[8] <= w61[8];
w62[9] <= w61[9];
w62[10] <= w61[10];
w62[11] <= w61[11];
w62[12] <= w61[12];
w62[13] <= w61[13];
w62[14] <= w61[14];
w62[15] <= w61[15];

a63 <= d62;
d63 <= c62;
c63 <= b62;
b63 <= b62 + (((a62 + (c62 ^ (b62 | (~d62))) + 'h2ad7d2bb + w62[(7 * 62) % 16]) << 15) | ((a62 + (c62 ^ (b62 | (~d62))) + 'h2ad7d2bb + w62[(7 * 62) % 16]) >> (32 - 15)));
w63[0] <= w62[0];
w63[1] <= w62[1];
w63[2] <= w62[2];
w63[3] <= w62[3];
w63[4] <= w62[4];
w63[5] <= w62[5];
w63[6] <= w62[6];
w63[7] <= w62[7];
w63[8] <= w62[8];
w63[9] <= w62[9];
w63[10] <= w62[10];
w63[11] <= w62[11];
w63[12] <= w62[12];
w63[13] <= w62[13];
w63[14] <= w62[14];
w63[15] <= w62[15];

a64 <= d63;
d64 <= c63;
c64 <= b63;
b64 <= b63 + (((a63 + (c63 ^ (b63 | (~d63))) + 'heb86d391 + w63[(7 * 63) % 16]) << 21) | ((a63 + (c63 ^ (b63 | (~d63))) + 'heb86d391 + w63[(7 * 63) % 16]) >> (32 - 21)));
		  
    end
endmodule



