`timescale 1ns / 1ns

module Md5CoreTest;

reg clk, reset, test_all;
wire [31:0] a, b, c, d;
reg [31:0] count = 0;
reg [511:0] chunk;

Md5Core m (
	.clk(clk), 
	.wb(chunk), 
	.a0('h67452301), 
	.b0('hefcdab89), 
	.c0('h98badcfe), 
	.d0('h10325476), 
	.a64(a), 
	.b64(b), 
	.c64(c), 
	.d64(d)
);


BytesToDWord converter(
  .byte0('hde),
  .byte1('had),
  .byte2('hbe),
  .byte3('hef)
);

initial
  begin
    clk = 0;
    forever #10 clk = !clk;
  end
  
initial
  begin
    reset = 0;
    #5 reset = 1;
    #4 reset = 0;
  end
  
initial
    $monitor($stime,, reset,, clk,,, count);    
    
`define TestCase(__number, __passed, __a, __b, __c, __d, __chunk)                           \
reg __passed;                                                                               \
always @(posedge clk)                                                                       \
  begin                                                                                     \
    if (count == __number)                                                                  \
      begin                                                                                 \
        chunk <= __chunk;                                                                   \
      end                                                                                   \
                                                                                            \
    if (count == __number + 65) __passed <= a == __a && b == __b && c == __c && d == __d;   \
  end                                                                                       \

`TestCase(
  0, 
  test0,
  'h35a8f271,
  'h39f4f1f4,
  'ha75fb5d4,
  'h4fba4572,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000)

`TestCase(
  1, 
  test1,
  'h7c9b108f,
  'hd07a467c,
  'h7352ebc5,
  'ha395f402,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100001)

`TestCase(
  2, 
  test2,
  'h89f035b0,
  'h376153aa,
  'h786deec9,
  'he4b6a605,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100010)

`TestCase(
  3, 
  test3,
  'h0eb78800,
  'h31c66081,
  'ha7618869,
  'h0d21345a,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100011)

`TestCase(
  4, 
  test4,
  'h6f38c6c2,
  'h22e7d460,
  'he70eab58,
  'hadda1dc0,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100100)

`TestCase(
  5, 
  test5,
  'h5db4ab0a,
  'h9ed72cd2,
  'h526b3edc,
  'h59960c96,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100101)

`TestCase(
  6, 
  test6,
  'h10bfdc6b,
  'hd2cd45cb,
  'h2cef75ac,
  'h3a7d9ea5,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100110)

`TestCase(
  7, 
  test7,
  'h23866d34,
  'hf7ec1067,
  'hb980578e,
  'hb940e343,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100111)

`TestCase(
  8, 
  test8,
  'h0bbfa183,
  'h3ee1a0b8,
  'h8ff6cad6,
  'he488f3c8,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000101000)

`TestCase(
  9, 
  test9,
  'h3b924e92,
  'hb0b9035a,
  'hd88cce0c,
  'h4cf3496d,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000101001)

`TestCase(
  10, 
  test10,
  'h7c956632,
  'hc0ac03d8,
  'hd7d3bf4e,
  'hb5daa1e1,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000101010)

`TestCase(
  11, 
  test11,
  'hbe2d8e25,
  'ha32d7b2d,
  'h3de4a73a,
  'h50ad5698,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000101011)

`TestCase(
  12, 
  test12,
  'ha81aa8bf,
  'hc3cc7846,
  'h3b41e4db,
  'hebecaaa9,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000101100)

`TestCase(
  13, 
  test13,
  'h55194a32,
  'h5e858acb,
  'hcab3f463,
  'h1771a867,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000101101)

`TestCase(
  14, 
  test14,
  'h48ac354f,
  'h4f95dcfa,
  'h1ef2bf62,
  'h8daa20e4,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000101110)

`TestCase(
  15, 
  test15,
  'h0f884365,
  'h5688be70,
  'h05289ea0,
  'hc994b7ff,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000101111)

`TestCase(
  16, 
  test16,
  'h1cdbaace,
  'hff982a0c,
  'h61250a68,
  'hca323383,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000110000)

`TestCase(
  17, 
  test17,
  'hd0fda7c3,
  'h92560e17,
  'h0195ef0f,
  'h8b5220f9,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000110001)

`TestCase(
  18, 
  test18,
  'h262cfbc7,
  'h7361a114,
  'hf0c42971,
  'h1c53c056,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000110010)

`TestCase(
  19, 
  test19,
  'h1783a8eb,
  'h0f14b0c2,
  'h40d4532a,
  'he388537c,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000110011)

`TestCase(
  20, 
  test20,
  'h12b15ca7,
  'h2e1a4819,
  'he2eba493,
  'h1bdfedff,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000110100)

`TestCase(
  21, 
  test21,
  'h17f6b7e3,
  'h55562332,
  'h6d709ad9,
  'hc4e64efe,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000110101)

`TestCase(
  22, 
  test22,
  'hb4c45615,
  'hbf41dcd1,
  'h702bd871,
  'hcc805d08,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000110110)

`TestCase(
  23, 
  test23,
  'hf89ef18e,
  'h8a493f45,
  'h4523595c,
  'h32f395d5,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000110111)

`TestCase(
  24, 
  test24,
  'h2eb3cdc8,
  'ha1dded72,
  'h3765185b,
  'h5cf129b3,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000111000)

`TestCase(
  25, 
  test25,
  'h6747a144,
  'hcdb181a5,
  'hb9413dec,
  'h167b7251,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000111001)

`TestCase(
  26, 
  test26,
  'ha8a41784,
  'h5b64a57a,
  'h7ceb61d9,
  'h0742f470,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000111010)

`TestCase(
  27, 
  test27,
  'h7472c99d,
  'h909f25d0,
  'h38b79f43,
  'he1c9a06b,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000111011)

`TestCase(
  28, 
  test28,
  'h110b2751,
  'h90cbcc98,
  'hf3d0cb23,
  'hc8aa745e,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000111100)

`TestCase(
  29, 
  test29,
  'hf5f9c942,
  'h7aa2c365,
  'h66b499f9,
  'h10f4fd74,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000111101)

`TestCase(
  30, 
  test30,
  'h3948bccd,
  'h64edbacb,
  'h1aada572,
  'h7f754050,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000111110)

`TestCase(
  31, 
  test31,
  'h0b3622d0,
  'h4a65503a,
  'hc1579428,
  'h4d78ea79,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000111111)

`TestCase(
  32, 
  test32,
  'h2e8d6b50,
  'hfbbec79c,
  'hb0e1e7dc,
  'hc376ba70,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000)

`TestCase(
  33, 
  test33,
  'h091da27e,
  'hb841fc5e,
  'h1e7a7c1c,
  'h198c57b8,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000001)

`TestCase(
  34, 
  test34,
  'h11913b9c,
  'hdaeeac75,
  'hfc852463,
  'h6183a604,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000010)

`TestCase(
  35, 
  test35,
  'hd0b33e0c,
  'h51500183,
  'hb4fda331,
  'h46dfe99e,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000011)

`TestCase(
  36, 
  test36,
  'hf3a200f5,
  'hcb94636a,
  'h5cb260d9,
  'ha584b73f,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000100)

`TestCase(
  37, 
  test37,
  'ha55b1b39,
  'h3c658a73,
  'h512b19ef,
  'hca61da2d,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000101)

`TestCase(
  38, 
  test38,
  'h2cd2e37f,
  'h6f6379a7,
  'h8693c188,
  'h01ddf293,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000110)

`TestCase(
  39, 
  test39,
  'h68e3acde,
  'hb69b99ea,
  'he901b6a8,
  'haf308a1e,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000111)

`TestCase(
  40, 
  test40,
  'ha8b0b6c0,
  'h2a8cd6fd,
  'h8c312525,
  'h863f6cd3,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001001000)

`TestCase(
  41, 
  test41,
  'h11f152dc,
  'ha0f1b7c2,
  'he718f2ee,
  'h6f4ac025,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001001001)

`TestCase(
  42, 
  test42,
  'ha31221fe,
  'ha173d741,
  'h23f4934a,
  'h75a8b7bb,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001001010)

`TestCase(
  43, 
  test43,
  'h3a81d0a4,
  'hadb55792,
  'h1be4d248,
  'h788f42c6,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001001011)

`TestCase(
  44, 
  test44,
  'h5c68e9d1,
  'hff50df2b,
  'h31f96f18,
  'h76f3660b,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001001100)

`TestCase(
  45, 
  test45,
  'h13d74668,
  'h7e011853,
  'hc858ad5f,
  'h9bd1d97c,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001001101)

`TestCase(
  46, 
  test46,
  'h14eb798c,
  'hb3f7482e,
  'h80ea452a,
  'h9a9c7cac,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001001110)

`TestCase(
  47, 
  test47,
  'h0fdc63f0,
  'habae17ca,
  'hf7d2b8a1,
  'h5e1db3ec,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001001111)

`TestCase(
  48, 
  test48,
  'h74599f43,
  'h825a8e87,
  'h73f23cf7,
  'h9aa7bb24,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001010000)

`TestCase(
  49, 
  test49,
  'h621f72ef,
  'h1db7ab41,
  'h98f8f94e,
  'hdde80028,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001010001)

`TestCase(
  50, 
  test50,
  'h6d8ebee0,
  'h8e44c77c,
  'h738e03a0,
  'hc650be39,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001010010)

`TestCase(
  51, 
  test51,
  'h7553995c,
  'h17d9d840,
  'h944de02a,
  'h5e21f2a4,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001010011)

`TestCase(
  52, 
  test52,
  'h259cc9b8,
  'h0b2d5f0c,
  'h6220326d,
  'hc2ffa2d9,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001010100)

`TestCase(
  53, 
  test53,
  'hf8fe3e4b,
  'hb0f2e851,
  'hba73d543,
  'hdb1f8d07,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001010101)

`TestCase(
  54, 
  test54,
  'ha310e351,
  'h1860bea7,
  'h39c4665c,
  'hbe2596e2,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001010110)

`TestCase(
  55, 
  test55,
  'h077bc660,
  'h608cfd20,
  'h46dec78a,
  'h66a003ee,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001010111)

`TestCase(
  56, 
  test56,
  'h5155ef01,
  'h2a4f5ad8,
  'h959e4f07,
  'h738171b7,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001011000)

`TestCase(
  57, 
  test57,
  'hac7fab56,
  'h977eb5f2,
  'h0a6971cd,
  'hd070af5a,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001011001)

`TestCase(
  58, 
  test58,
  'h2ea09f20,
  'h11a41ca8,
  'ha38ff658,
  'hc54f57ba,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001011010)

`TestCase(
  59, 
  test59,
  'hbed23180,
  'h0528caf6,
  'h86ebc762,
  'hcb2d6327,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001011011)

`TestCase(
  60, 
  test60,
  'h8152b027,
  'h73ea5aea,
  'h751d6121,
  'he003390f,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001011100)

`TestCase(
  61, 
  test61,
  'h0ed29a0e,
  'hd5550258,
  'h3ac5939c,
  'hcba22ae6,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001011101)

`TestCase(
  62, 
  test62,
  'h96e5477d,
  'h8a3872cc,
  'h37401d77,
  'h71a751d1,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001011110)

`TestCase(
  63, 
  test63,
  'h193627b0,
  'h65f32dd0,
  'hced76f97,
  'h21ce91d6,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001011111)

`TestCase(
  64, 
  test64,
  'ha351023d,
  'habf92ff0,
  'h54196f69,
  'h51fa52f1,
  'b00000000000000000000000000000000000000000000000000000000010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000110010001101100011100100110111101110111001000000110111101101100011011000110010101001000)

`TestCase(
  65, 
  test65,
  'h35e1d885,
  'h955e6190,
  'hf38c03f8,
  'h0ff85076,
  'b00000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000010110010001101100011100100110111101110111001000000110111101101100011011000110010101001000)

`TestCase(
  66, 
  test66,
  'h3637ed9d,
  'h92e87fae,
  'h9c62fb6d,
  'hc5e74fcc,
  'b00000000000000000000000000000000000000000000000000000001010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001100111011011110110010000100000011110010111101001100001011011000010000001100101011010000111010000100000011100100110010101110110011011110010000001110011011100000110110101110101011010100010000001111000011011110110011000100000011011100111011101101111011100100110001000100000011010110110001101101001011101010111000100100000011001010110100001010100)

`TestCase(
  67, 
  test67,
  'h5ac4b6e3,
  'h2d2e2507,
  'h15448ba2,
  'hc098ce69,
  'b00000000000000000000000000000000000000000000000000000001011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010111001100111011011110110010000100000011110010111101001100001011011000010000001100101011010000111010000100000011100100110010101110110011011110010000001110011011100000110110101110101011010100010000001111000011011110110011000100000011011100111011101101111011100100110001000100000011010110110001101101001011101010111000100100000011001010110100001010100)

`TestCase(
  68, 
  test68,
  'hfb44bc89,
  'h5b68a719,
  'ha7550760,
  'hdb9d42ca,
  'b00000000000000000000000000000000000000000000000000000000010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000110100001100011011101000110100101100101010011000010000001101110011010000110111101001010)
  
    
always @(posedge clk)
  begin
    count <= count + 1;
  end 
  
always @(posedge test68)
  test_all <= test0&test1&test2&test3&test4&test5&test6&test7&test8&test9&test10&test11&test12&test13&test14&test15&test16&test17&test18&test19&test20&test21&test22&test23&test24&test25&test26&test27&test28&test29&test30&test31&test32&test33&test34&test35&test36&test37&test38&test39&test40&test41&test42&test43&test44&test45&test46&test47&test48&test49&test50&test51&test52&test53&test54&test55&test56&test57&test58&test59&test60&test61&test62&test63&test64&test65&test66&test67&test68;
    
endmodule  

 

